module m41 (parameter N = 4) (input [N-1:0] A, B, C, D 
output [1:0] SEL, [N-1:0] OUT);


endmodule