module equality_comparator(input [N-1:0] A, B, output OUT);

assign OUT = (A == B);

endmodule