module full_adder_tb;
logic a = 0;
logic b = 0;
logic cin = 0;

wire cout, sum;

endmodule